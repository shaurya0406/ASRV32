`timescale 1ns/1ps
`default_nettype none

`include "asrv32_header.vh"

/* ALU Module & Ports Declaration*/
module asrv32_alu
    (
        /* Inputs */
        input wire i_clk,i_rst_n,               // Input Clock & Active Low Reset
        // ! We have clock enable now | input wire i_alu_en,                    // Enable Signal indicating the ALU stage (EXE stage) is currently active
        
        /* From Decoder */
        input wire[31:0] i_pc_idex,
        input wire[4:0] i_rs1_addr_idex,
        input wire[4:0] i_rs2_addr_idex,
        input wire[4:0] i_rd_addr_idex,
        input wire[31:0] i_imm_idex,                 // Immediate value generated by Decoder from previous stage (ID)
        input wire[2:0] i_funct3_idex,
        input wire[`OPCODE_WIDTH-1:0] i_opcode_idex, // Instruction Opcode Type from previous stage (ID)
        input wire[`ALU_WIDTH-1:0] i_alu_op_idex,    // ALU operation type from previous stage (ID)
        input wire[`EXCEPTION_WIDTH-1:0] i_exception_idex,
        
        /* From BaseReg (DECODE Stage) */
        input wire[31:0] i_rs1_data,            // Data read from the first source register.
        input wire[31:0] i_rs2_data,            // Data read from the second source register.
        
        // ! PC Value
        // ! now we get PC from pipeline prev stage (ID) | input wire[31:0] i_pc,  // PC value from FETCH Stage (IF)

        /* Memory */
        output reg[31:0] o_alu_result_exmem,     // Result of arithmetic operation by ALU
        output reg[31:0] o_rs2_data_exmem,       // Data to be stored to memory is always rs2
        
        /* CSR */
        output reg[4:0] o_rs1_addr_excsr,
        output reg[31:0] o_rs1_data_excsr,
        output reg[11:0] o_imm_excsr, // ! 12 bits only
        output reg[`EXCEPTION_WIDTH-1:0] o_exception_excsr,

        /* Common to Memory & CSR */
        output reg[2:0] o_funct3_exmemcsr,
        output reg[`OPCODE_WIDTH-1:0] o_opcode_exmemcsr,

        /* PC Control */
        output reg[31:0] o_pc_exmem,    // pc register in pipeline
        output reg[31:0] o_next_pc,     // new pc value
        output reg o_change_pc,         // high if PC needs to jump

        /* BaseReg Control */
        output reg o_wr_rd, //write rd to the base reg if enabled
        input wire[4:0] i_rd_addr, //address for destination register (from previous stage)
        output reg[4:0] o_rd_addr, //address for destination register
        output reg[31:0] o_rd_data, //value to be written back to destination register
        output reg o_rd_valid, //high if o_rd_data is valid (not load nor csr instruction)
        
        /* Pipeline Control */
        output reg o_stall_from_alu, //prepare to stall next stage(memory-access stage) for load/store instruction
        input wire i_ce, // Global clk enable for pipeline stalling of this stage
        output reg o_ce, // Global clk enable for pipeline stalling of next stage
        input wire i_stall, // informs this stage to stall
        input wire i_force_stall, // ! force this stage to stall in case of hazard
        output reg o_stall, // informs pipeline to stall
        input wire i_flush, // flush this stage
        output reg o_flush // flush previous stages
    );

// ! will move this to testbench
// /* For Testbench */
//     initial begin
//         o_alu_result = 0;
//     end

/* Intermediate Register Declaration: */
    reg[31:0] y_d;  // Store ALU Result
    reg[31:0] a;    // Store Operand 1
    reg[31:0] b;    // Store Operand 2
    reg[31:0] rd_data_d; // Next value to be written back to destination register
    reg wr_rd_d;    // Write rd to basereg if enabled
    reg rd_valid_d; // High if rd is valid (neither load nor csr instruction)
    reg[31:0] a_pc; 
    wire[31:0] sum;

/* Internal Parallel Wires for less resource utilisation */
    wire alu_add    = i_alu_op_idex[`ADD];
    wire alu_sub    = i_alu_op_idex[`SUB];
    wire alu_slt    = i_alu_op_idex[`SLT];
    wire alu_sltu   = i_alu_op_idex[`SLTU];
    wire alu_xor    = i_alu_op_idex[`XOR];
    wire alu_or     = i_alu_op_idex[`OR];
    wire alu_and    = i_alu_op_idex[`AND];
    wire alu_sll    = i_alu_op_idex[`SLL];
    wire alu_srl    = i_alu_op_idex[`SRL];
    wire alu_sra    = i_alu_op_idex[`SRA];
    wire alu_eq     = i_alu_op_idex[`EQ];
    wire alu_neq    = i_alu_op_idex[`NEQ];
    wire alu_ge     = i_alu_op_idex[`GE];
    wire alu_geu    = i_alu_op_idex[`GEU];

    wire opcode_rtype = i_opcode_idex[`RTYPE];
    wire opcode_itype = i_opcode_idex[`ITYPE];
    wire opcode_load = i_opcode_idex[`LOAD];
    wire opcode_store = i_opcode_idex[`STORE];
    wire opcode_branch = i_opcode_idex[`BRANCH];
    wire opcode_jal = i_opcode_idex[`JAL];
    wire opcode_jalr = i_opcode_idex[`JALR];
    wire opcode_lui = i_opcode_idex[`LUI];
    wire opcode_auipc = i_opcode_idex[`AUIPC];
    wire opcode_system = i_opcode_idex[`SYSTEM];
    wire opcode_fence = i_opcode_idex[`FENCE];

/* Stall Logic for this stage (EX) */
    wire stall_bit  = o_stall || i_stall;

/* ALU Arithmetic Combinational Logic (Blocking Code): */
    always @* begin  
        y_d = 0;                        // Default value of intermediate register y_d
        a = (opcode_jal || opcode_auipc)    ? i_pc_idex :i_rs1_data;    // a can either be pc or rs1
        b = (opcode_rtype || opcode_branch) ? i_rs2_data:i_imm_idex;    // b can either be rs2 or imm 

        if(alu_add) y_d = a + b;        // Addition
        if(alu_sub) y_d = a - b;        // Subtraction
        if(alu_slt || alu_sltu) begin   // Set if less than
            y_d = {31'b0, (a < b)};                // Less than comparison
            if(alu_slt) y_d = (a[31] ^ b[31])? {31'b0,a[31]}:y_d;   // Consider sign bit for signed comparison
        end 
        if(alu_xor) y_d = a ^ b;        // Bitwise XOR
        if(alu_or)  y_d = a | b;        // Bitwise OR
        if(alu_and) y_d = a & b;        // Bitwise AND
        if(alu_sll) y_d = a << b[4:0];  // Shift left logical
        if(alu_srl) y_d = a >> b[4:0];  // Shift right logical
        if(alu_sra) y_d = $signed(a) >>> b[4:0]; // Shift right arithmetic
        if(alu_eq || alu_neq) begin     // Equality check
            y_d = {31'b0,(a == b)};               // Check if equal
            if(alu_neq) y_d = {31'b0,!y_d[0]};     // Invert result for not equal
        end
        if(alu_ge || alu_geu) begin     // Greater than or equal check
            y_d = {31'b0,(a >= b)};               // Check if greater than or equal
            if(alu_ge) y_d = (a[31] ^ b[31])? {31'b0, b[31]}:y_d;    // Consider sign bit for signed comparison
        end
    end

/* Determine o_rd_data and Next PC Value */
    always @* begin
        o_flush = i_flush; //flush this stage along with the previous stages
        rd_data_d = 0;
        rd_valid_d = 0;
        o_change_pc = 0;
        o_next_pc = 0;
        wr_rd_d = 0;
        a_pc = i_pc_idex;
        if(!i_flush) begin
            if(opcode_rtype || opcode_itype) rd_data_d = y_d;
            if(opcode_branch && y_d[0]) begin
                    o_next_pc = sum; //branch iff value of ALU is 1(true)
                    o_change_pc = i_ce; //change PC when ce of this stage is high (o_change_pc is valid)
                    o_flush = i_ce;
            end
            if(opcode_jal || opcode_jalr) begin
                if(opcode_jalr) a_pc = i_rs1_data;
                o_next_pc = sum; //jump to new PC
                o_change_pc = i_ce; //change PC when ce of this stage is high (o_change_pc is valid)
                o_flush = i_ce;
                rd_data_d = i_pc_idex + 4; //register the next pc value to destination register
            end 
        end
        if(opcode_lui) rd_data_d = i_imm_idex;
        if(opcode_auipc) rd_data_d = sum;

        if(opcode_branch || opcode_store || (opcode_system && i_funct3_idex == 0) || opcode_fence ) wr_rd_d = 0; //i_funct3_idex==0 are the non-csr system instructions 
        else wr_rd_d = 1; //always write to the destination reg except when instruction is BRANCH or STORE or SYSTEM(except CSR system instruction)  

        if(opcode_load || (opcode_system && i_funct3_idex!=0)) rd_valid_d = 0;  //value of o_rd_data for load and CSR write is not yet available at this stage
        else rd_valid_d = 1;

        //stall logic (stall when upper stages are stalled, when forced to stall, or when needs to flush previous stages but are still stalled)
        o_stall = (i_stall || i_force_stall) && !i_flush; //stall when alu needs wait time
    end
        
    assign sum = a_pc + i_imm_idex; //share adder for all addition operation for less resource utilization

/* Register the ALU Output */
    always @(posedge i_clk, negedge i_rst_n) begin
        if(!i_rst_n) begin
            o_exception_excsr   <= 0;
            o_ce                <= 0;
            o_stall_from_alu    <= 0;
        end
        else begin
           if(i_ce && !stall_bit) begin //update register only if this stage is enabled
                o_opcode_exmemcsr   <= i_opcode_idex;
                o_exception_excsr   <= i_exception_idex;
                o_alu_result_exmem  <= y_d; 
                o_rs1_addr_excsr    <= i_rs1_addr_idex;
                o_rs1_data_excsr    <= i_rs1_data;
                o_rs2_data_exmem    <= i_rs2_data;
                o_rd_addr           <= i_rd_addr_idex;
                o_imm_excsr         <= i_imm_idex[11:0];
                o_funct3_exmemcsr   <= i_funct3_idex;
                o_rd_data           <= rd_data_d;
                o_rd_valid          <= rd_valid_d;
                o_wr_rd             <= wr_rd_d;
                o_stall_from_alu    <= i_opcode_idex[`STORE] || i_opcode_idex[`LOAD]; //stall next stage(memory-access stage) when need to store/load since accessing data memory always takes more than 1 cycle
                o_pc_exmem          <= i_pc_idex;
            end
            if(i_flush && !stall_bit) begin //flush this stage so clock-enable of next stage is disabled at next clock cycle
                o_ce <= 0;
            end
            else if(!stall_bit) begin //clock-enable will change only when not stalled
                o_ce <= i_ce;
            end
            else if(stall_bit && !i_stall) o_ce <= 0; //if this stage is stalled but next stage is not, disable clock enable of next stage at next clock cycle (pipeline bubble) 
        end
    end 

endmodule